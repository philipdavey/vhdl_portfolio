-- ====================================================================
-- File Name     : <insert_file_name>
-- Author        : Philip Davey
-- Design Folder : <insert_design_folder>
-- Date          : <insert_date>
-- Rtl/Sim/Pkg   : <insert>
-- --------------------------------------------------------------------
-- HDL           : <insert>
-- --------------------------------------------------------------------
-- Description   :
--               :
--               :
--               :
--               :
-- ====================================================================