PACKAGE aes_pkg IS

    TYPE S_BOX_ARRAY IS ARRAY (15 DOWNTO 0) OF STD_LOGIC_VECTOR(31 DOWNTO 0);
    CONSTANT S_BOX

END PACKAGE aes_pkg;

PACKAGE BODY aes_pkg IS

END PACKAGE BODY aes_pkg;
